module top_module (
    output out);
    
    out=0; //it takes as decimal by default

endmodule
